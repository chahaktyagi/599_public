module stage_ID_EX (
    input           ID__stage_ID_EX_regwrite,
    input           ID__stage_ID_EX_memtoreg,
    input           ID__stage_ID_EX_memread,
    input           ID__stage_ID_EX_memwrite,
    input           ID__stage_ID_EX_alusrc,
    input   [1:0]   ID__stage_ID_EX_aluop,
    input           ID__stage_ID_EX_regdst,
    input           ID__stage_ID_EX_sys_en,
    input   [31:0]  ID__stage_ID_EX_rs_data,
    input   [31:0]  ID__stage_ID_EX_rt_data,
    input   [4:0]   ID__stage_ID_EX_rs_id,
    input   [4:0]   ID__stage_ID_EX_rt_id,
    input   [4:0]   ID__stage_ID_EX_rd_id,
    input   [31:0]  ID__stage_ID_EX_sign_ext,
    input   [2:0]   ID__stage_ID_EX_funct3,
    output          stage_ID_EX__EX_regwrite,
    output          stage_ID_EX__EX_memtoreg,
    output          stage_ID_EX__EX_memread,
    output          stage_ID_EX__EX_memwrite,
    output          stage_ID_EX__EX_alusrc,
    output   [1:0]  stage_ID_EX__EX_aluop,
    output          stage_ID_EX__EX_regdst,
    output          stage_ID_EX__EX_sys_en,
    output   [31:0] stage_ID_EX__EX_rs_data,
    output   [31:0] stage_ID_EX__EX_rt_data,
    output   [4:0]  stage_ID_EX__EX_rs_id,
    output   [4:0]  stage_ID_EX__EX_rt_id,
    output   [4:0]  stage_ID_EX__EX_rd_id,
    output   [31:0] stage_ID_EX__EX_sign_ext,
    output   [2:0]  stage_ID_EX__EX_funct3
);
endmodule